library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ALU is
    port (
        alu_A : in std_logic_vector(15 downto 0);
        alu_B : in std_logic_vector(15 downto 0);
        instr : in integer;
        alu_C : out std_logic_vector(15 downto 0);
        C, Z  : out std_logic
    );
end entity ALU;

architecture rtl of ALU is

    function perform_addition(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
        variable C_par       : std_logic := '0';
        variable G, P        : std_logic;
    begin
        add_instance: for i in 0 to 15 loop
            G := A(i) and B(i);
            P := A(i) xor B(i);
            temp_result(i) := P xor C_par;
            C_par := G or (P and C_par);
        end loop add_instance;						
        return temp_result;
    end function;

     function perform_4bit_addition(A, B : std_logic_vector(3 downto 0); Cin: std_logic) return std_logic_vector is
        variable temp_result : std_logic_vector(4 downto 0);
        variable C_par       : std_logic := Cin;
        variable G, P        : std_logic;
    begin
        add_instance: for i in 0 to 3 loop
            G := A(i) and B(i);
            P := A(i) xor B(i);
            temp_result(i) := P xor C_par;
            C_par := G or (P and C_par);
        end loop add_instance;
	    temp_result(4) := C_par;
        return temp_result;
    end function;

    function perform_subtraction(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
        variable C_par       : std_logic := '1';
        variable G, P        : std_logic;
    begin
        sub_instance: for i in 0 to 15 loop
            G := A(i) and (not B(i));
            P := A(i) xor (not B(i));
            temp_result(i) := P xor C_par;
            C_par := G or (P and C_par);
        end loop sub_instance;						  
        return temp_result;
    end function;    

    function perform_multiplication(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
        variable product     : std_logic_vector(7 downto 0) := "00000000";
	variable AB0,AB1,AB2,AB3,t1a,t2a,t3a : std_logic_vector(3 downto 0);
	variable t1,t2,t3: std_logic_vector(5 downto 0);
    begin
	k1: for i in 0 to 3 loop:
	begin
		AB0(i) <= A(i) and B(0);
		AB1(i) <= A(i) and B(1);
		AB2(i) <= A(i) and B(2);
		AB3(i) <= A(i) and B(3);
	end loop k1;

	
	t1a(2 downto 0) := AB0(3 downto 1);
	t1a(3) := '0';
	t1 := perform_4bit_addition(t1a,AB1,'0');
	t2a(2 downto 0) := t1(3 downto 1);
	t2a(3) := '0';
	t2 := perform_4bit_addition(t2a,AB2,t1a(4));
	t3a(2 downto 0) := t2(3 downto 1);
	t3a(3) := '0';
	t3 := perform_4bit_addition(t3a,AB3,t2a(4));
	temp_result(0) := AB0(0);
	temp_result(1) := t1(0);
	temp_result(2) := t2(0);
	temp_result(7 downto 3) := t3;
        return temp_result;
    end function;    

    function perform_and(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
    begin
        and_instance: for i in 0 to 15 loop
            temp_result(i) := A(i) and B(i);
        end loop and_instance;
        return temp_result;
    end function;    

    function perform_or(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
    begin
        or_instance: for i in 0 to 15 loop
            temp_result(i) := A(i) or B(i);
        end loop or_instance;
        return temp_result;
    end function;    

    function perform_imp(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
    begin
        imp_instance: for i in 0 to 15 loop
            temp_result(i) := (not A(i)) or B(i);
        end loop imp_instance;
        return temp_result;
    end function;    

    function perform_LLI(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
        variable A_par       : std_logic_vector(8 downto 0) := A(8 downto 0);
        variable B_par       : std_logic_vector(6 downto 0) := B(6 downto 0);
    begin
        temp_result := A_par & B_par;
        return temp_result;
    end function;    

    function perform_LHI(A, B : std_logic_vector(15 downto 0)) return std_logic_vector is
        variable temp_result : std_logic_vector(15 downto 0);
        variable A_par       : std_logic_vector(8 downto 0) := A(8 downto 0);
        variable B_par       : std_logic_vector(6 downto 0) := B(6 downto 0);
    begin
        temp_result := B_par & A_par;
        return temp_result;
    end function;    

    function carry_flag(A, B: std_logic_vector(15 downto 0); M: std_logic) return std_logic is
        variable result : std_logic := M;
        variable G, P   : std_logic;
    begin 
        add_instance: for i in 0 to 15 loop 
            G := A(i) and B(i);
            P := A(i) xor B(i);
            result := G or (P and result);
        end loop add_instance;
        return result;
    end function;    

    function z_flag(A, B: std_logic_vector(15 downto 0)) return std_logic is
        variable result : std_logic;
        variable subtraction : std_logic_vector(15 downto 0) := perform_subtraction(A, B);
    begin
        z_instance: if subtraction = "0000000000000000" generate
                        result := '1';
                    else 
                        result := '0'; 
                    end generate z_instance;
    
        return result;
    end function;    
  
begin 
    with instr select
        alu_C <= perform_addition(alu_A, alu_B)       when 1,
                 perform_subtraction (alu_A, alu_B)   when 2,
                 perform_multiplication(alu_A, alu_B) when 3,
                 perform_and(alu_A, alu_B)            when 4,
                 perform_or(alu_A, alu_B)	          when 5,
                 perform_imp(alu_A, alu_B)	          when 6,
                 perfomr_LHI(alu_A, alu_B)	          when 7,
	             perfomr_LLI(alu_A, alu_B)	          when 8;

    with instr select 
        C <= carry_flag(alu_A, alu_B, '0') when 1,
             carry_flag(alu_A, alu_B, '1') when 2,
             '0' when others;
             
    with instr select 
        Z <= z_flag(alu_A, alu_B) when 2,
             '0' when others;

end architecture;
